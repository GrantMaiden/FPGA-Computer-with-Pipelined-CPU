/*
memory functions as a static RAM, with 2K (2048) x 16-bit memory locations.
From an external view, memory functionally has 1K (1024) x 32-bit memory locations.
This means that addresses entered into this module are assumed to range from 0 to 1023.

memory supports RW operations, executing these operations using a 32-bit I/O port.

To operate memory, clear chip_select to select the device and enable R/W operations. 
Reading: Clear output enable, enter address into MAR, set RW
Writing: Set output enable, enter address and write data in MDR, and clear RW

Note: Signals in memory propagate after delay (example: when reading, it will take
a propagation delay after entering an address to display memory's data).

Note: Reset operation is NOT supported in memory module, as it is too costly
to wipe the memory module.
*/
module memory #(parameter DEPTH=2048, parameter FILE="sample.txt")
               (clk, reset, data, address, out_en, chip_s, RW);
   input  logic clk, reset;     // Clock, Reset signals
	inout  [31:0] data;          // Bidirectional 32-bit I/O port
	// 11-bit address input- see Note.
	input  logic [9:0] address;
	// Output enable: 1 to write to data, 0 to read from data
   input  logic out_en;
	// Chip select: 1 to disable R/W, 0 to enable R/W
	input  logic chip_s;
   // Read/Write: 1 to read, 0 to write to memory
	// Assume write takes place on posedge of RW (if RW is strobed for one cycle)
	// Note: If write is held low for more than one cycle, data is simply written until
	// one cycle after RW goes high.
	input  logic RW;
	
	// Initial Logic
	// 
	initial begin
		$readmemh(FILE, stored_memory);
	end
	
	
	// Memory Address Registers: Adjacent addresses
	logic  [10:0] MAR1, MAR2;
	assign MAR1 = (address * 11'd2);
	assign MAR2 = ((address * 11'd2) + 11'd1);
	
	// Memory Data Registers: higher bits and lower bits
	logic  [15:0] MDRHigh, MDRLow;

	// 16-bit values with a parameterized depth
	logic [15:0] stored_memory [(DEPTH-1):0];
	
	always_ff @(posedge clk) begin
		if (!RW /*&& !out_en*/ && !chip_s) begin            // Write to memory
			stored_memory[MAR1] <= data[31:16];
			stored_memory[MAR2] <=  data[15:0];
		end
	end
	
	// Combinational Logic
	// Output enable behavior:
	// If 1, IO port gets high Z (Write)
	// If 0, IO port gets data_out (Read)
	/*assign data[31:16] = (!out_en && !chip_s && RW) ? MDRHigh : 16'bZ;
	assign  data[15:0] = (!out_en && !chip_s && RW) ?  MDRLow : 16'bZ;*/
	
	assign data = (!out_en && !chip_s && RW) ? {MDRHigh, MDRLow} : 32'bz;
	
	// Sequential Logic
	always_ff @(posedge clk) begin
		if (RW && !out_en /*&& !chip_s*/) begin            // Read from memory
			MDRHigh <= stored_memory[MAR1];
			MDRLow  <= stored_memory[MAR2];
		end
	end
	
endmodule

// Tester Module
module memory_testbench();
	logic clk, reset;     // Clock, Reset signals
	wire  [31:0] data;    // Bidirectional 32-bit I/O port
	logic [9:0] address; // !!! Note: Takes 0-1023 (10 bits max)
   logic out_en;
	logic chip_s;
	logic RW;
	
	// Local value to feed IO port when writing
	logic [31:0] data1;
	
	memory dut (clk, reset, data, address, out_en, chip_s, RW);
	
	// Note: when ACCESSING memory, output enable logic is inverted
	// (depending which way you define it)
	// ...
	// Need to add chip select, all those other signals...
//	assign data = (out_en) ? data1 : 16'bz;
	assign data[31:0] = (out_en) ? data1 : 32'bz;
	
	// Set up the clock.
	parameter CLOCK_PERIOD=100;
	initial begin
		clk <= 0;
		forever #(CLOCK_PERIOD/2) clk <= ~clk;
	end
	
	// Set up the inputs to the design. Each line is a clock cycle.
	// Test... set direction to pass data in
	// Then clear direction to read data
	initial begin
								  @(posedge clk);
	chip_s <= 0; 	        @(posedge clk);
								  @(posedge clk);
	RW <= 1;               @(posedge clk);
								  @(posedge clk);
	out_en <= 1; address <= 10'b1111111111; data1 <= 65555; @(posedge clk);
								  @(posedge clk);
								  @(posedge clk);
	RW <= 0;               @(posedge clk);
	RW <= 1;               @(posedge clk);
								  @(posedge clk);
								  @(posedge clk);
	address <= 10'b01; data1 <= 25050; @(posedge clk);
								  @(posedge clk);
	RW <= 0;               @(posedge clk);
	RW <= 1;               @(posedge clk);
	address <= 10'b01000; data1 <= 2; @(posedge clk);
								  @(posedge clk);
	RW <= 0;               @(posedge clk);
	RW <= 1;               @(posedge clk);
								  @(posedge clk);
								  @(posedge clk);
	out_en <= 0; address <= 11'b010; @(posedge clk);
								  @(posedge clk);
	address <= 10'b01;     @(posedge clk);
	address <= 10'b01000;  @(posedge clk);
////	out_en <= 1; address <= 11'b00; data1 <= {16{1'b1}}; data2 <= {16{1'b1}}; @(posedge clk);
//	out_en <= 1; address <= 11'b00; data1 <= {16{1'b1}}; data2 <= {16{1'b0}}; @(posedge clk);
//								  @(posedge clk);
//								  @(posedge clk);
//	RW <= 0;               @(posedge clk);
//	RW <= 1;               @(posedge clk);
//								  @(posedge clk);
//								  @(posedge clk);
//	address <= 11'b01; data1 <= {16{1'b0}}; data2 <= {16{1'b0}}; @(posedge clk);
//								  @(posedge clk);
//	RW <= 0;               @(posedge clk);
//	RW <= 1;               @(posedge clk);
//	address <= 11'b01000; data1 <= 16'b0000111100001111; data2 <= 16'b0000111100001111; @(posedge clk);
//								  @(posedge clk);
//	RW <= 0;               @(posedge clk);
//	RW <= 1;               @(posedge clk);
//								  @(posedge clk);
//								  @(posedge clk);
//	out_en <= 0; address <= 11'b010; @(posedge clk);
//								  @(posedge clk);
//	address <= 11'b01;     @(posedge clk);
//	address <= 11'b01000;  @(posedge clk);
								  @(posedge clk);
								  @(posedge clk);
								  @(posedge clk);
								  @(posedge clk);
//	out_en <= 1; address <= 4'b0111; data1 <= 4'b0000; @(posedge clk);
//	RW <= 0;               @(posedge clk);
//	RW <= 1;               @(posedge clk);
//	out_en <= 0;           @(posedge clk);
//	address <= 4'b0110;    @(posedge clk);
//								  @(posedge clk);
//	address <= 4'b0000;    @(posedge clk);
								  @(posedge clk);
								  @(posedge clk);
	$stop; // End the simulation.
	end
endmodule
